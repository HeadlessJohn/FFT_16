`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////

module TB_16();
    reg clk;
    reg rst;
    reg signed [15:0] data_0, data_1, data_2, data_3, data_4, data_5, data_6, data_7;
    reg signed [15:0] data_8, data_9, data_10, data_11, data_12, data_13, data_14, data_15;

    wire signed [15:0] o_f0_r, o_f1_r, o_f2_r, o_f3_r, o_f4_r, o_f5_r, o_f6_r, o_f7_r;
    wire signed [15:0] o_f8_r, o_f9_r, o_f10_r, o_f11_r, o_f12_r, o_f13_r, o_f14_r, o_f15_r;

    wire signed [15:0] o_f0_i, o_f1_i, o_f2_i, o_f3_i, o_f4_i, o_f5_i, o_f6_i, o_f7_i;
    wire signed [15:0] o_f8_i, o_f9_i, o_f10_i, o_f11_i, o_f12_i, o_f13_i, o_f14_i, o_f15_i;

    // wire [22:0] f0, f1, f2, f3, f4, f5, f6, f7;
    initial begin
        clk = 0;
        rst = 1;
        #20
        rst = 0;
        forever #10 clk = ~clk; // 20MHz
    end

    initial begin
        
         

        #20    
        // sin 1wave
        data_0 =  0      *(127);// + 127;
        data_1 =  0.3826 *(127);// + 127;
        data_2 =  0.7071 *(127);// + 127;
        data_3 =  0.9238 *(127);// + 127;
        data_4 =  1      *(127);// + 127;
        data_5 =  0.9238 *(127);// + 127;
        data_6 =  0.7071 *(127);// + 127;
        data_7 =  0.3826 *(127);// + 127;
        data_8 =  0      *(127);// + 127;
        data_9 =  -0.3826*(127);// + 127;
        data_10 = -0.7071*(127);// + 127;
        data_11 = -0.9238*(127);// + 127;
        data_12 = -1     *(127);// + 127;
        data_13 = -0.9238*(127);// + 127;
        data_14 = -0.7071*(127);// + 127;
        data_15 = -0.3826*(127);// + 127;
    
        #20
        // sin 2wave
        data_0  = 0       *(127);// + 127; 
        data_1  = 0.7071  *(127);// + 127;      
        data_2  = 1       *(127);// + 127;    
        data_3  = 0.7071  *(127);// + 127;      
        data_4  = 0       *(127);// + 127;     
        data_5  = -0.7071 *(127);// + 127;  
        data_6  = -1      *(127);// + 127;    
        data_7  = -0.7071 *(127);// + 127;   
        data_8  = 0       *(127);// + 127;   
        data_9  = 0.7071  *(127);// + 127;    
        data_10 = 1       *(127);// + 127;    
        data_11 = 0.7071  *(127);// + 127;  
        data_12 = 0       *(127);// + 127;   
        data_13 = -0.7071 *(127);// + 127;  
        data_14 = -1      *(127);// + 127;  
        data_15 = -0.7071 *(127);// + 127;   
        
        #20
        // sin 3wave
        data_0  = 0 *(127);// + 127; 
        data_1  = 0.9238 *(127);// + 127;      
        data_2  = 0.7071 *(127);// + 127;    
        data_3  = -0.3826 *(127);// + 127;      
        data_4  = -1 *(127);// + 127;     
        data_5  = -0.3826 *(127);// + 127;  
        data_6  = 0.7071 *(127);// + 127;    
        data_7  = 0.9238 *(127);// + 127;   
        data_8  = 0 *(127);// + 127;   
        data_9  = -0.9238 *(127);// + 127;    
        data_10 = -0.7071 *(127);// + 127;    
        data_11 = 0.3826 *(127);// + 127;  
        data_12 = 1 *(127);// + 127;   
        data_13 = 0.3826 *(127);// + 127;  
        data_14 = -0.7071 *(127);// + 127;  
        data_15 = -0.9238 *(127);// + 127;   

        #20
        // sin 4wave
        data_0  = 0 *(127);// + 127; 
        data_1  = 1 *(127);// + 127;      
        data_2  = 0 *(127);// + 127;    
        data_3  = -1 *(127);// + 127;      
        data_4  = 0 *(127);// + 127;     
        data_5  = 1 *(127);// + 127;  
        data_6  = 0 *(127);// + 127;    
        data_7  = -1 *(127);// + 127;   
        data_8  = 0 *(127);// + 127;   
        data_9  = 1 *(127);// + 127;    
        data_10 = 0 *(127);// + 127;    
        data_11 = -1 *(127);// + 127;  
        data_12 = 0 *(127);// + 127;   
        data_13 = 1 *(127);// + 127;  
        data_14 = 0 *(127);// + 127;  
        data_15 = -1 *(127);// + 127;   

        #20
        // sin 5wave
        data_0  = 0 *(127);// + 127; 
        data_1  = 0.9238 *(127);// + 127;      
        data_2  = -0.7071 *(127);// + 127;    
        data_3  = -0.3826 *(127);// + 127;      
        data_4  = 1 *(127);// + 127;     
        data_5  = -0.3826 *(127);// + 127;  
        data_6  = -0.7071 *(127);// + 127;    
        data_7  = 0.9238 *(127);// + 127;   
        data_8  = 0 *(127);// + 127;   
        data_9  = -0.9238 *(127);// + 127;    
        data_10 = 0.7071 *(127);// + 127;    
        data_11 = 0.3826 *(127);// + 127;  
        data_12 = -1 *(127);// + 127;   
        data_13 = 0.3826 *(127);// + 127;  
        data_14 = 0.7071 *(127);// + 127;  
        data_15 = -0.9238 *(127);// + 127;   

        #20
        // sin 6wave
        data_0 =  0       *(127);// + 127;
        data_1 =  0.7071 *(127);// + 127;
        data_2 =  -1 *(127);// + 127;
        data_3 =  0.7071 *(127);// + 127;
        data_4 =  0 *(127);// + 127;
        data_5 =  -0.7071 *(127);// + 127;
        data_6 =  1 *(127);// + 127;
        data_7 =  -0.7071 *(127);// + 127;
        data_8 =  0 *(127);// + 127;
        data_9 =  0.7071 *(127);// + 127;
        data_10 = -1 *(127);// + 127;
        data_11 = 0.7071 *(127);// + 127;
        data_12 = 0 *(127);// + 127;
        data_13 = -0.7071 *(127);// + 127;
        data_14 = 1 *(127);// + 127;
        data_15 = -0.7071 *(127);// + 127;
        
        #20
        // sin 7wave
        data_0  = 0 *(127);// + 127;  
        data_1  = 0.3826 *(127);// + 127; 
        data_2  = -0.7071 *(127);// + 127;      
        data_3  = 0.9238 *(127);// + 127;    
        data_4  = -1 *(127);// + 127;      
        data_5  = 0.9238 *(127);// + 127;     
        data_6  = -0.7071 *(127);// + 127;  
        data_7  = 0.3826 *(127);// + 127;    
        data_8  = 0 *(127);// + 127;   
        data_9  = -0.3826 *(127);// + 127;   
        data_10 = 0.7071 *(127);// + 127;    
        data_11 = -0.9238 *(127);// + 127;    
        data_12 = 1 *(127);// + 127;  
        data_13 = -0.9238 *(127);// + 127;   
        data_14 = 0.7071 *(127);// + 127;  
        data_15 = -0.3826 *(127);// + 127;  

        #20
        // cos 1wave
        data_0 =  1      *(127);// + 127;
        data_1 =  0.9238 *(127);// + 127;
        data_2 =  0.7071 *(127);// + 127;
        data_3 =  0.3826 *(127);// + 127;
        data_4 =  0      *(127);// + 127;
        data_5 =  -0.3826*(127);// + 127;
        data_6  = -0.7071*(127);// + 127;
        data_7  = -0.9238*(127);// + 127;
        data_8  = -1     *(127);// + 127;
        data_9  = -0.9238*(127);// + 127;
        data_10 = -0.7071*(127);// + 127;
        data_11 = -0.3826*(127);// + 127;
        data_12 =  0      *(127);// + 127;
        data_13 =  0.3826 *(127);// + 127;
        data_14 =  0.7071 *(127);// + 127;
        data_15 =  0.9238 *(127);// + 127

        #20
        // cos 2wave
        data_0  = 1       *(127);// + 127;    
        data_1  = 0.7071  *(127);// + 127;      
        data_2  = 0       *(127);// + 127;     
        data_3  = -0.7071 *(127);// + 127;  
        data_4  = -1      *(127);// + 127;    
        data_5  = -0.7071 *(127);// + 127;   
        data_6  = 0       *(127);// + 127;   
        data_7  = 0.7071  *(127);// + 127;    
        data_8  = 1       *(127);// + 127;    
        data_9  = 0.7071  *(127);// + 127;  
        data_10 = 0       *(127);// + 127;   
        data_11 = -0.7071 *(127);// + 127;  
        data_12 = -1      *(127);// + 127;  
        data_13 = -0.7071 *(127);// + 127;   
        data_14 = 0       *(127);// + 127; 
        data_15 = 0.7071  *(127);// + 127;    

        #20
        // cos 3wave
        data_0  = 1 *(127);// + 127;   
        data_1  = 0.3826 *(127);// + 127;  
        data_2  = -0.7071 *(127);// + 127;  
        data_3  = -0.9238 *(127);// + 127;     
        data_4  = 0 *(127);// + 127; 
        data_5  = 0.9238 *(127);// + 127;      
        data_6  = 0.7071 *(127);// + 127;    
        data_7  = -0.3826 *(127);// + 127;      
        data_8  = -1 *(127);// + 127;     
        data_9  = -0.3826 *(127);// + 127;  
        data_10 = 0.7071 *(127);// + 127;    
        data_11 = 0.9238 *(127);// + 127;   
        data_12 = 0 *(127);// + 127;   
        data_13 = -0.9238 *(127);// + 127;    
        data_14 = -0.7071 *(127);// + 127;    
        data_15 = 0.3826 *(127);// + 127;  

        #20
        // cos 4wave
        data_0  = 1 *(127);// + 127;      
        data_1  = 0 *(127);// + 127;    
        data_2  = -1 *(127);// + 127;      
        data_3  = 0 *(127);// + 127;     
        data_4  = 1 *(127);// + 127;  
        data_5  = 0 *(127);// + 127;    
        data_6  = -1 *(127);// + 127;   
        data_7  = 0 *(127);// + 127;   
        data_8  = 1 *(127);// + 127;    
        data_9  = 0 *(127);// + 127;    
        data_10 = -1 *(127);// + 127;  
        data_11 = 0 *(127);// + 127;   
        data_12 = 1 *(127);// + 127;  
        data_13 = 0 *(127);// + 127;  
        data_14 = -1 *(127);// + 127;   
        data_15 = 0 *(127);// + 127; 

        #20
        // cos 5wave
        data_0  = 1 *(127);// + 127;     
        data_1  = -0.3826 *(127);// + 127;  
        data_2  = -0.7071 *(127);// + 127;    
        data_3  = 0.9238 *(127);// + 127;   
        data_4  = 0 *(127);// + 127;   
        data_5  = -0.9238 *(127);// + 127;    
        data_6  = 0.7071 *(127);// + 127;    
        data_7  = 0.3826 *(127);// + 127;  
        data_8  = -1 *(127);// + 127;   
        data_9  = 0.3826 *(127);// + 127;  
        data_10 = 0.7071 *(127);// + 127;  
        data_11 = -0.9238 *(127);// + 127;   
        data_12 = 0 *(127);// + 127; 
        data_13 = 0.9238 *(127);// + 127;      
        data_14 = -0.7071 *(127);// + 127;    
        data_15 = -0.3826 *(127);// + 127;      

        #20
        // cos 6wave
        data_0  = 1 *(127);// + 127;
        data_1  = -0.7071 *(127);// + 127;
        data_2 =  0       *(127);// + 127;
        data_3 =  0.7071 *(127);// + 127;
        data_4 =  -1 *(127);// + 127;
        data_5 =  0.7071 *(127);// + 127;
        data_6 =  0 *(127);// + 127;
        data_7 =  -0.7071 *(127);// + 127;
        data_8 =  1 *(127);// + 127;
        data_9 =  -0.7071 *(127);// + 127;
        data_10=  0 *(127);// + 127;
        data_11=  0.7071 *(127);// + 127;
        data_12 = -1 *(127);// + 127;
        data_13 = 0.7071 *(127);// + 127;
        data_14 = 0 *(127);// + 127;
        data_15 = -0.7071 *(127);// + 127;
        
        #20
        // cos 7wave
        data_0  = 1 *(127);// + 127;  
        data_1  = -0.9238 *(127);// + 127;   
        data_2  = 0.7071 *(127);// + 127;  
        data_3  = -0.3826 *(127);// + 127;  
        data_4  = 0 *(127);// + 127;  
        data_5  = 0.3826 *(127);// + 127; 
        data_6  = -0.7071 *(127);// + 127;      
        data_7  = 0.9238 *(127);// + 127;    
        data_8  = -1 *(127);// + 127;      
        data_9  = 0.9238 *(127);// + 127;     
        data_10 = -0.7071 *(127);// + 127;  
        data_11 = 0.3826 *(127);// + 127;    
        data_12 = 0 *(127);// + 127;   
        data_13 = -0.3826 *(127);// + 127;   
        data_14 = 0.7071 *(127);// + 127;    
        data_15 = -0.9238 *(127);// + 127;    

        #20
        // cos 8wave
        data_0  = 1 *(127); 
        data_1  = -1*(127);
        data_2  = 1 *(127); 
        data_3  = -1*(127);
        data_4  = 1 *(127); 
        data_5  = -1*(127);
        data_6  = 1 *(127); 
        data_7  = -1*(127);
        data_8  = 1 *(127); 
        data_9  = -1*(127);
        data_10 = 1 *(127); 
        data_11 = -1*(127);
        data_12 = 1 *(127); 
        data_13 = -1*(127);
        data_14 = 1 *(127); 
        data_15 = -1*(127);

        #20
        // dc
        data_0  = 1*(127); 
        data_1  = 1*(127);
        data_2  = 1*(127); 
        data_3  = 1*(127);
        data_4  = 1*(127); 
        data_5  = 1*(127);
        data_6  = 1*(127); 
        data_7  = 1*(127);
        data_8  = 1*(127); 
        data_9  = 1*(127);
        data_10 = 1*(127); 
        data_11 = 1*(127);
        data_12 = 1*(127); 
        data_13 = 1*(127);
        data_14 = 1*(127); 
        data_15 = 1*(127);
        // #10
        // 3sin3x + sinx
        // data_0  = 0; 
        // data_1  = 100;
        // data_2  = 90; 
        // data_3  = -7;
        // data_4  = -64; 
        // data_5  = -7;
        // data_6  = 90; 
        // data_7  = 100;
        // data_8  = 0; 
        // data_9  = -100;
        // data_10 = -90; 
        // data_11 = 7;
        // data_12 = 64; 
        // data_13 = 7;
        // data_14 = -90; 
        // data_15 = -100;

        #10
        // 2cos2x + sin3x
        // data_0  =   84;
        // data_1  =   98;
        // data_2  =   29;
        // data_3  =  -76;
        // data_4  =  -127;
        // data_5  =  -76;
        // data_6  =   29;
        // data_7  =   98;
        // data_8  =   84;
        // data_9  =   20;
        // data_10 =  -29;
        // data_11 =  -43;
        // data_12 =  -42;
        // data_13 =  -43;
        // data_14 =  -29;
        // data_15 =   20;

        #10
        // sinx + 2sin2x + 3sin3x
        // data_0  =     0 + 30;
        // data_1  =    96 + 30;
        // data_2  =   102 + 30;
        // data_3  =    25 + 30;
        // data_4  =   -42 + 30;
        // data_5  =   -34 + 30;
        // data_6  =    17 + 30;
        // data_7  =    36 + 30;
        // data_8  =     0 + 30;
        // data_9  =   -36 + 30;
        // data_10 =   -17 + 30;
        // data_11 =    34 + 30;
        // data_12 =    42 + 30;
        // data_13 =   -25 + 30;
        // data_14 =  -102 + 30;
        // data_15 =   -96 + 30;

        #10
        // 3cosx + 2cos2x + cos3x + sin3x
        // data_0  =   84 + 40;
        // data_1  =   77 + 40;
        // data_2  =   29 + 40;
        // data_3  =  -22 + 40;
        // data_4  =  -42 + 40;
        // data_5  =  -28 + 40;
        // data_6  =   -9 + 40;
        // data_7  =  -11 + 40;
        // data_8  =  -28 + 40;
        // data_9  =  -37 + 40;
        // data_10 =  -29 + 40;
        // data_11 =  -17 + 40;
        // data_12 =  -14 + 40;
        // data_13 =  -11 + 40;
        // data_14 =    9 + 40;
        // data_15 =   51 + 40;

        // #20
        // // dc
        // data_0  = 8'd1;
        // data_1  = 8'd1;
        // data_2  = 8'd1;
        // data_3  = 8'd1;
        // data_4  = 8'd1;
        // data_5  = 8'd1;
        // data_6  = 8'd1;
        // data_7  = 8'd1;
        // data_8  = 8'd1;
        // data_9  = 8'd1;
        // data_10 = 8'd1;
        // data_11 = 8'd1;
        // data_12 = 8'd1;
        // data_13 = 8'd1;
        // data_14 = 8'd1;
        // data_15 = 8'd1;

        #80 $stop;
        #10
        // sin 8wave
        data_0  = 0;
        data_1  = 0;
        data_2  = 0;
        data_3  = 0;
        data_4  = 0;
        data_5  = 0;
        data_6  = 0;
        data_7  = 0;
        data_8  = 0;
        data_9  = 0;
        data_10 = 0;
        data_11 = 0;
        data_12 = 0;
        data_13 = 0;
        data_14 = 0;
        data_15 = 0;



        // sin 9wave
        // data_0 =  0       *(127);// + 127;
        // data_1 =  -0.3826 *(127);// + 127;
        // data_2 =  0.7071  *(127);// + 127;
        // data_3 =  -0.9238 *(127);// + 127;
        // data_4 =  1       *(127);// + 127;
        // data_5 =  -0.9238 *(127);// + 127;
        // data_6 =  0.7071  *(127);// + 127;
        // data_7 =  -0.3826 *(127);// + 127;
        // data_8 =  0       *(127);// + 127;
        // data_9 =  0.3826  *(127);// + 127;
        // data_10 = -0.7071 *(127);// + 127;
        // data_11 =  0.9238 *(127);// + 127;
        // data_12 =  -1     *(127);// + 127;
        // data_13 =  0.9238 *(127);// + 127;
        // data_14 =  -0.7071*(127);// + 127;
        // data_15 =  0.3826 *(127);// + 127;

        // cosin 2wave
        // data_0  =  0      *(127);// + 127;
        // data_1  =  -0.7071*(127);// + 127;
        // data_2  =  -1     *(127);// + 127;
        // data_3  =  -0.7071*(127);// + 127;
        // data_4  =  0      *(127);// + 127;
        // data_5  =  0.7071 *(127);// + 127;
        // data_6   =  1      *(127);// + 127;
        // data_7   =  0.7071 *(127);// + 127;
        // data_8   =  0      *(127);// + 127;
        // data_9   =  -0.7071*(127);// + 127;
        // data_10  =  -1     *(127);// + 127;
        // data_11  =  -0.7071*(127);// + 127;
        // data_12 =  0      *(127);// + 127;
        // data_13 =  0.7071 *(127);// + 127;
        // data_14 =  1      *(127);// + 127;
        // data_15 =  0.7071 *(127);// + 127;



        // square
        // data_0  = 8'd255;
        // data_1  = 8'd0;
        // data_2  = 8'd255;
        // data_3  = 8'd0;
        // data_4  = 8'd255;
        // data_5  = 8'd0;
        // data_6  = 8'd255;
        // data_7  = 8'd0;
        // data_8  = 8'd255;
        // data_9  = 8'd0;
        // data_10 = 8'd255;
        // data_11 = 8'd0;
        // data_12 = 8'd255;
        // data_13 = 8'd0;
        // data_14 = 8'd255;
        // data_15 = 8'd0;

    end
    
    FFT_16 DUT_01(
        .clk(clk),
        .rst(rst),
        .data_0(data_0), 
        .data_1(data_1), 
        .data_2(data_2), 
        .data_3(data_3), 
        .data_4(data_4), 
        .data_5(data_5), 
        .data_6(data_6), 
        .data_7(data_7),
        .data_8(data_8),
        .data_9(data_9),
        .data_10(data_10),
        .data_11(data_11),
        .data_12(data_12),
        .data_13(data_13),
        .data_14(data_14),
        .data_15(data_15),
        .o_f0_r(o_f0_r), 
        .o_f0_i(o_f0_i), 
        .o_f1_r(o_f1_r), 
        .o_f1_i(o_f1_i), 
        .o_f2_r(o_f2_r), 
        .o_f2_i(o_f2_i), 
        .o_f3_r(o_f3_r), 
        .o_f3_i(o_f3_i), 
        .o_f4_r(o_f4_r), 
        .o_f4_i(o_f4_i), 
        .o_f5_r(o_f5_r), 
        .o_f5_i(o_f5_i), 
        .o_f6_r(o_f6_r),
        .o_f6_i(o_f6_i),
        .o_f7_r(o_f7_r),
        .o_f7_i(o_f7_i),
        .o_f8_r(o_f8_r), 
        .o_f8_i(o_f8_i), 
        .o_f9_r(o_f9_r), 
        .o_f9_i(o_f9_i), 
        .o_f10_r(o_f10_r), 
        .o_f10_i(o_f10_i), 
        .o_f11_r(o_f11_r), 
        .o_f11_i(o_f11_i), 
        .o_f12_r(o_f12_r), 
        .o_f12_i(o_f12_i), 
        .o_f13_r(o_f13_r), 
        .o_f13_i(o_f13_i), 
        .o_f14_r(o_f14_r),
        .o_f14_i(o_f14_i),
        .o_f15_r(o_f15_r),
        .o_f15_i(o_f15_i)
    );

    // abs_sum abs(
    //     .f0_r(o_f0_r),
    //     .f0_i(o_f0_i),
    //     .f1_r(o_f1_r),
    //     .f1_i(o_f1_i),
    //     .f2_r(o_f2_r),
    //     .f2_i(o_f2_i),
    //     .f3_r(o_f3_r),
    //     .f3_i(o_f3_i),
    //     .f4_r(o_f4_r),
    //     .f4_i(o_f4_i),
    //     .f5_r(o_f5_r),
    //     .f5_i(o_f5_i),
    //     .f6_r(o_f6_r),
    //     .f6_i(o_f6_i),
    //     .f7_r(o_f7_r),
    //     .f7_i(o_f7_i),
    //     .f0(f0), 
    //     .f1(f1), 
    //     .f2(f2), 
    //     .f3(f3), 
    //     .f4(f4), 
    //     .f5(f5), 
    //     .f6(f6), 
    //     .f7(f7)
    // );

endmodule


module TB_FFT_16_total();
    reg [15:0] data_in;
    
    reg [19:0] sampling_period;
    reg [3:0] read_addr;

    wire [15:0] data_r;
    wire [15:0] data_i;

    wire sampling_signal;
    wire [3:0] write_addr;

    reg clk, rst;

   initial begin
        clk = 0;
        rst = 1;
        #10
        rst = 0;
        data_in = 0;
        sampling_period = 50;
        read_addr = 0;
        forever #10 clk = ~clk; // 20MHz
    end

    initial begin
        repeat(100) begin
            #20
            data_in = 10;
            #20
            data_in = 30;
            #20
            data_in = 60;
            #20
            data_in = 100;
            #20
            data_in = 60;
            #20
            data_in = 30;
            #20
            data_in = 10;
            #20
            data_in = 0;
            read_addr = read_addr + 1;
        end
        $stop;
    end

	sampling_clk samp_inst(
		.clk(clk),
		.rst(rst),
		.sampling_period(sampling_period), // 1_048_575 clocks
		.sampling_signal(sampling_signal)
    );

	addr_cnt addr_inst(
		.clk(clk),
		.rst(rst),
		.clk_in(sampling_signal),
		.addr(write_addr)
    );

	TOP top_inst(
		.clk(clk),
		.rst(rst),
		.data_in(data_in),
		.write_addr(write_addr),
		.we(1),
		.read_addr(read_addr),
		.re(1),
		.data_r(data_r),
		.data_i(data_i)
    );
endmodule